// Copyright (C) 2016  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel MegaCore Function License Agreement, or other 
// applicable license agreement, including, without limitation, 
// that your use is for the sole purpose of programming logic 
// devices manufactured by Intel and sold by Intel or its 
// authorized distributors.  Please refer to the applicable 
// agreement for further details.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 16.1.1 Build 200 11/30/2016 SJ Lite Edition"
// CREATED		"Mon Feb 13 18:12:47 2017"

module project02_la(
	D,
	S
);


input wire	[3:0] D;
output wire	[6:0] S;

wire	test;
wire	SYNTHESIZED_WIRE_0;
wire	SYNTHESIZED_WIRE_1;
wire	SYNTHESIZED_WIRE_78;
wire	SYNTHESIZED_WIRE_79;
wire	SYNTHESIZED_WIRE_80;
wire	SYNTHESIZED_WIRE_81;
wire	SYNTHESIZED_WIRE_9;
wire	SYNTHESIZED_WIRE_10;
wire	SYNTHESIZED_WIRE_11;
wire	SYNTHESIZED_WIRE_12;
wire	SYNTHESIZED_WIRE_19;
wire	SYNTHESIZED_WIRE_20;
wire	SYNTHESIZED_WIRE_21;
wire	SYNTHESIZED_WIRE_22;
wire	SYNTHESIZED_WIRE_23;
wire	SYNTHESIZED_WIRE_24;
wire	SYNTHESIZED_WIRE_32;
wire	SYNTHESIZED_WIRE_33;
wire	SYNTHESIZED_WIRE_34;
wire	SYNTHESIZED_WIRE_35;
wire	SYNTHESIZED_WIRE_36;
wire	SYNTHESIZED_WIRE_37;
wire	SYNTHESIZED_WIRE_41;
wire	SYNTHESIZED_WIRE_42;
wire	SYNTHESIZED_WIRE_43;
wire	SYNTHESIZED_WIRE_44;
wire	SYNTHESIZED_WIRE_54;
wire	SYNTHESIZED_WIRE_55;
wire	SYNTHESIZED_WIRE_56;
wire	SYNTHESIZED_WIRE_57;
wire	SYNTHESIZED_WIRE_58;
wire	SYNTHESIZED_WIRE_59;
wire	SYNTHESIZED_WIRE_63;
wire	SYNTHESIZED_WIRE_64;
wire	SYNTHESIZED_WIRE_65;
wire	SYNTHESIZED_WIRE_68;
wire	SYNTHESIZED_WIRE_69;
wire	SYNTHESIZED_WIRE_74;
wire	SYNTHESIZED_WIRE_75;
wire	SYNTHESIZED_WIRE_76;
wire	SYNTHESIZED_WIRE_77;




assign	SYNTHESIZED_WIRE_79 =  ~D[3];

assign	SYNTHESIZED_WIRE_81 =  ~D[2];

assign	S[0] = SYNTHESIZED_WIRE_0 | SYNTHESIZED_WIRE_1;

assign	SYNTHESIZED_WIRE_11 = D[0] & SYNTHESIZED_WIRE_78 & D[3];

assign	SYNTHESIZED_WIRE_10 = D[0] & test & SYNTHESIZED_WIRE_79;

assign	SYNTHESIZED_WIRE_12 = SYNTHESIZED_WIRE_80 & SYNTHESIZED_WIRE_78 & SYNTHESIZED_WIRE_79;

assign	SYNTHESIZED_WIRE_9 = SYNTHESIZED_WIRE_80 & SYNTHESIZED_WIRE_81;

assign	SYNTHESIZED_WIRE_68 = SYNTHESIZED_WIRE_9 | SYNTHESIZED_WIRE_10 | SYNTHESIZED_WIRE_11 | SYNTHESIZED_WIRE_12;

assign	SYNTHESIZED_WIRE_21 = SYNTHESIZED_WIRE_78 & SYNTHESIZED_WIRE_79;

assign	SYNTHESIZED_WIRE_20 = D[0] & SYNTHESIZED_WIRE_79;

assign	SYNTHESIZED_WIRE_22 = D[0] & SYNTHESIZED_WIRE_78;

assign	SYNTHESIZED_WIRE_19 = D[2] & SYNTHESIZED_WIRE_79;

assign	SYNTHESIZED_WIRE_78 =  ~test;

assign	SYNTHESIZED_WIRE_24 = SYNTHESIZED_WIRE_81 & D[3];

assign	SYNTHESIZED_WIRE_23 = SYNTHESIZED_WIRE_19 | SYNTHESIZED_WIRE_20 | SYNTHESIZED_WIRE_21 | SYNTHESIZED_WIRE_22;

assign	S[2] = SYNTHESIZED_WIRE_23 | SYNTHESIZED_WIRE_24;

assign	SYNTHESIZED_WIRE_34 = SYNTHESIZED_WIRE_78 & D[3];

assign	SYNTHESIZED_WIRE_33 = SYNTHESIZED_WIRE_80 & SYNTHESIZED_WIRE_81 & SYNTHESIZED_WIRE_79;

assign	SYNTHESIZED_WIRE_35 = D[0] & test & SYNTHESIZED_WIRE_81;

assign	SYNTHESIZED_WIRE_32 = D[0] & SYNTHESIZED_WIRE_78 & D[2];

assign	SYNTHESIZED_WIRE_37 = SYNTHESIZED_WIRE_80 & test & D[2];

assign	SYNTHESIZED_WIRE_36 = SYNTHESIZED_WIRE_32 | SYNTHESIZED_WIRE_33 | SYNTHESIZED_WIRE_34 | SYNTHESIZED_WIRE_35;

assign	S[3] = SYNTHESIZED_WIRE_36 | SYNTHESIZED_WIRE_37;

assign	SYNTHESIZED_WIRE_80 =  ~D[0];

assign	SYNTHESIZED_WIRE_43 = SYNTHESIZED_WIRE_80 & SYNTHESIZED_WIRE_81;

assign	SYNTHESIZED_WIRE_42 = SYNTHESIZED_WIRE_80 & test;

assign	SYNTHESIZED_WIRE_44 = test & D[3];

assign	SYNTHESIZED_WIRE_41 = D[2] & D[3];

assign	S[4] = SYNTHESIZED_WIRE_41 | SYNTHESIZED_WIRE_42 | SYNTHESIZED_WIRE_43 | SYNTHESIZED_WIRE_44;

assign	SYNTHESIZED_WIRE_56 = SYNTHESIZED_WIRE_81 & D[3];

assign	SYNTHESIZED_WIRE_55 = test & D[3];

assign	SYNTHESIZED_WIRE_57 = SYNTHESIZED_WIRE_80 & SYNTHESIZED_WIRE_78 & SYNTHESIZED_WIRE_79;

assign	SYNTHESIZED_WIRE_54 = SYNTHESIZED_WIRE_78 & D[2] & SYNTHESIZED_WIRE_79;

assign	SYNTHESIZED_WIRE_59 = SYNTHESIZED_WIRE_80 & test & D[2];

assign	SYNTHESIZED_WIRE_76 = SYNTHESIZED_WIRE_81 & SYNTHESIZED_WIRE_80;

assign	SYNTHESIZED_WIRE_58 = SYNTHESIZED_WIRE_54 | SYNTHESIZED_WIRE_55 | SYNTHESIZED_WIRE_56 | SYNTHESIZED_WIRE_57;

assign	S[5] = SYNTHESIZED_WIRE_58 | SYNTHESIZED_WIRE_59;

assign	SYNTHESIZED_WIRE_63 = SYNTHESIZED_WIRE_78 & D[2];

assign	SYNTHESIZED_WIRE_65 = SYNTHESIZED_WIRE_80 & test;

assign	SYNTHESIZED_WIRE_64 = test & SYNTHESIZED_WIRE_81;

assign	S[6] = SYNTHESIZED_WIRE_63 | SYNTHESIZED_WIRE_64 | D[3] | SYNTHESIZED_WIRE_65;

assign	SYNTHESIZED_WIRE_69 = SYNTHESIZED_WIRE_81 & SYNTHESIZED_WIRE_79;

assign	S[1] = SYNTHESIZED_WIRE_68 | SYNTHESIZED_WIRE_69;

assign	SYNTHESIZED_WIRE_75 = test & SYNTHESIZED_WIRE_79;

assign	SYNTHESIZED_WIRE_77 = D[2] & test;

assign	SYNTHESIZED_WIRE_74 = D[0] & D[2] & SYNTHESIZED_WIRE_79;

assign	SYNTHESIZED_WIRE_1 = SYNTHESIZED_WIRE_78 & SYNTHESIZED_WIRE_81 & D[3];

assign	SYNTHESIZED_WIRE_0 = SYNTHESIZED_WIRE_74 | SYNTHESIZED_WIRE_75 | SYNTHESIZED_WIRE_76 | SYNTHESIZED_WIRE_77;

assign	test = D[1];

endmodule
